module image_rom(
   input wire [4:0] row,
   output [479:0] rgb);
	
reg [479:0] data; 

always @*
      case (row)
         0: data <= 479'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff; 
			1: data <= 479'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
			2: data <= {96'hffffffffffffffffffffffff, {8'h0, 4'hf}, 12'h000, 240'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff, 12'h000, {8'h0, 4'hf}, 96'hffffffffffffffffffffffff};
			3: data <= {84'hfffffffffffffffffffff, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {8'h0, 4'hf}, 12'h000, 204'hfffffffffffffffffffffffffffffffffffffffffffffffffff, 12'h000, {8'h0, 4'hf}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, 84'hfffffffffffffffffffff};
			4: data <= {84'hfffffffffffffffffffff, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {8'h0, 4'hf}, 12'h000, 96'hffffffffffffffffffffffff, 12'h000, 12'hfff, 24'h000, 60'hfffffffffffffff, 12'h000, {8'h0, 4'hf}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, 84'hfffffffffffffffffffff};
			5: data <= {96'hffffffffffffffffffffffff, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {8'h0, 4'hf}, 12'h000, 72'hffffffffffffffffff, 12'h000, {8'h0, 4'hf}, 12'h000, {8'h0, 4'hf}, 12'h000, 48'hffffffffffff, 12'h000, {8'h0, 4'hf}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, 84'hfffffffffffffffffffff};
			6: data <= {84'hfffffffffffffffffffff, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {8'h0, 4'hf}, 12'h000, 48'hffffffffffff, 12'h000, 12'h000, {8'h0, 4'hf}, 12'h000, {8'h0, 4'hf}, 12'h000, 12'h000, 48'hffffffffffff, 12'h000, {8'h0, 4'hf}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, 84'hfffffffffffffffffffff};
			7: data <= {84'hfffffffffffffffffffff, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {8'h0, 4'hf}, 24'hffffff, 12'h000, 12'h000, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, 12'h000, 12'h000, 24'hffffff, {8'h0, 4'hf}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, 96'hffffffffffffffffffffffff};
			8: data <= {84'hfffffffffffffffffffff, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {8'h0, 4'hf}, 12'hfff, 12'h000, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, 12'h000, 12'hfff, {8'h0, 4'hf}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, 84'hfffffffffffffffffffff};
			9: data <= {84'hfffffffffffffffffffff, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {8'h0, 4'hf}, 12'h000, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, 12'h000, {8'h0, 4'hf}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, 84'hfffffffffffffffffffff};
			10: data <= {96'hffffffffffffffffffffffff, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, 12'h000, {4'h6, 4'hb, 4'hf}, 12'h000, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, 12'h000, {4'h6, 4'hb, 4'hf}, 12'h000, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, {4'hf, 4'hb, 4'hc}, 96'hffffffffffffffffffffffff};
			11: data <= {96'hffffffffffffffffffffffff, 12'h000, {4'hf, 4'hb, 4'hc}, 12'h000, {4'h6, 4'hb, 4'hf}, 36'h000000000, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, 36'h000000000, {4'h6, 4'hb, 4'hf}, 12'h000, {4'hf, 4'hb, 4'hc}, 12'h000, 96'hffffffffffffffffffffffff};
			12: data <= {108'hfffffffffffffffffffffffffff, {4'hf, 4'hb, 4'hc}, 12'h000, {4'h6, 4'hb, 4'hf}, 24'h000000, 12'hfff, 12'h000, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, 12'h000, 12'hfff, 24'h000000, {4'h6, 4'hb, 4'hf}, 12'h000, {4'hf, 4'hb, 4'hc}, 108'hfffffffffffffffffffffffffff};
			13: data <= {108'hfffffffffffffffffffffffffff, 24'h000000, {4'h6, 4'hb, 4'hf}, 48'h000000000000, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, 48'h000000000000, {4'h6, 4'hb, 4'hf}, 24'h000000, 108'hfffffffffffffffffffffffffff};
			14: data <= {120'hffffffffffffffffffffffffffffff, 12'h000, {4'h6, 4'hb, 4'hf}, 12'h000, 12'hfff, 24'h000000, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, 36'h000000000, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, 24'h000000, 12'hfff, 12'h000, {4'h6, 4'hb, 4'hf}, 12'h000, 120'hffffffffffffffffffffffffffffff};
			15: data <= {120'hffffffffffffffffffffffffffffff, 12'h000, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, 24'h000000, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, 60'h000000000000000, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, 24'h000000, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, 12'h000, 120'hffffffffffffffffffffffffffffff};
			16: data <= {120'hffffffffffffffffffffffffffffff, 12'h000, {8'h0, 4'hf}, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, 36'h000000000, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, 12'h000, 120'hffffffffffffffffffffffffffffff};
			17: data <= {132'hfffffffffffffffffffffffffffffffff, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, 132'hfffffffffffffffffffffffffffffffff};
			18: data <= {144'hffffffffffffffffffffffffffffffffffff, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, 144'hffffffffffffffffffffffffffffffffffff};
			19: data <= {192'hffffffffffffffffffffffffffffffffffffffffffffffff, 12'h000, {8'h0, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {8'h0, 4'hf}, 12'h000, 192'hffffffffffffffffffffffffffffffffffffffffffffffff}; 
			20: data <= {180'hfffffffffffffffffffffffffffffffffffffffffffff, 12'h000, {8'h0, 4'hf}, {8'h0, 4'hf}, 12'h000, {4'h6, 4'hb, 4'hf}, 12'h000, {8'h0, 4'hf}, {8'h0, 4'hf}, 12'h000, 180'hfffffffffffffffffffffffffffffffffffffffffffff};
			21: data <= {168'hffffffffffffffffffffffffffffffffffffffffff, 36'h000000000, {8'h0, 4'hf}, 12'h000, {4'h6, 4'hb, 4'hf}, 12'h000, {8'h0, 4'hf}, 36'h000000000, 168'hffffffffffffffffffffffffffffffffffffffffff};
			22: data <= {156'hfffffffffffffffffffffffffffffffffffffff, 12'h000, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, 24'h000000, {4'h6, 4'hb, 4'hf}, 24'h000000, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, 12'h000, 156'hfffffffffffffffffffffffffffffffffffffff};
			23: data <= {156'hfffffffffffffffffffffffffffffffffffffff, 36'h000000000, {8'h0, 4'hf}, 12'h000, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, 12'h000, {8'h0, 4'hf}, 36'h000000000, 156'hfffffffffffffffffffffffffffffffffffffff};
			24: data <= {156'hfffffffffffffffffffffffffffffffffffffff, 36'h000000000, {8'h0, 4'hf}, 12'h000, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, {4'h6, 4'hb, 4'hf}, 12'h000, {8'h0, 4'hf}, 36'h000000000, 156'hfffffffffffffffffffffffffffffffffffffff};
			25: data <= {156'hfffffffffffffffffffffffffffffffffffffff, 12'h000, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, 60'h000000000000000, {8'h0, 4'hf}, {8'h0, 4'hf}, {8'h0, 4'hf}, 12'h000, 156'hfffffffffffffffffffffffffffffffffffffff};
			26: data <= {168'hffffffffffffffffffffffffffffffffffffffffff, 36'h000000000, 60'hfffffffffffffff, 36'h000000000, 168'hffffffffffffffffffffffffffffffffffffffffff};
			27: data <= 479'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
			28: data <= 479'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
			29: data <= 479'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
			
 endcase  
 
assign rgb = data;
 
 endmodule