//https://github.com/bogini/Pong/blob/master/font_rom.v

module font_rom(
    input wire clk,
    input wire [10:0] addr,
    output reg [7:0] data_reg
   );
	
reg [7:0] data; 
reg [10:0] addr_reg; 

always @(posedge clk) 
      addr_reg <= addr;

always @*
      case (addr_reg)
			//code x00
         11'h000: data <= 8'b00000000; // 
         11'h001: data <= 8'b00000000; // 
         11'h002: data <= 8'b00000000; // 
         11'h003: data <= 8'b00000000; // 
         11'h004: data <= 8'b00000000; // 
         11'h005: data <= 8'b00000000; // 
         11'h006: data <= 8'b00000000; // 
         11'h007: data <= 8'b00000000; // 
         11'h008: data <= 8'b00000000; // 
         11'h009: data <= 8'b00000000; // 
         11'h00a: data <= 8'b00000000; // 
         11'h00b: data <= 8'b00000000; // 
         11'h00c: data <= 8'b00000000; // 
         11'h00d: data <= 8'b00000000; // 
         11'h00e: data <= 8'b00000000; // 
         11'h00f: data <= 8'b00000000; // 
			//code x2a
         11'h2a0: data <= 8'b00000000; // 
         11'h2a1: data <= 8'b00000000; // 
         11'h2a2: data <= 8'b00000000; // 
         11'h2a3: data <= 8'b00000000; // 
         11'h2a4: data <= 8'b00000000; // 
         11'h2a5: data <= 8'b01100110; //  **  **
         11'h2a6: data <= 8'b00111100; //   ****
         11'h2a7: data <= 8'b11111111; // ********
         11'h2a8: data <= 8'b00111100; //   ****
         11'h2a9: data <= 8'b01100110; //  **  **
         11'h2aa: data <= 8'b00000000; // 
         11'h2ab: data <= 8'b00000000; // 
         11'h2ac: data <= 8'b00000000; // 
         11'h2ad: data <= 8'b00000000; // 
         11'h2ae: data <= 8'b00000000; // 
         11'h2af: data <= 8'b00000000; // 	
			//code x2b
         11'h2b0: data <= 8'b00000000; // 
         11'h2b1: data <= 8'b00000000; // 
         11'h2b2: data <= 8'b00000000; // 
         11'h2b3: data <= 8'b00000000; // 
         11'h2b4: data <= 8'b00000000; // 
         11'h2b5: data <= 8'b00011000; //    **
         11'h2b6: data <= 8'b00011000; //    **
         11'h2b7: data <= 8'b01111110; //  ******
         11'h2b8: data <= 8'b00011000; //    **
         11'h2b9: data <= 8'b00011000; //    **
         11'h2ba: data <= 8'b00000000; // 
         11'h2bb: data <= 8'b00000000; // 
         11'h2bc: data <= 8'b00000000; // 
         11'h2bd: data <= 8'b00000000; // 
         11'h2be: data <= 8'b00000000; // 
         11'h2bf: data <= 8'b00000000; // 
			//code x2d
         11'h2d0: data <= 8'b00000000; // 
         11'h2d1: data <= 8'b00000000; // 
         11'h2d2: data <= 8'b00000000; // 
         11'h2d3: data <= 8'b00000000; // 
         11'h2d4: data <= 8'b00000000; // 
         11'h2d5: data <= 8'b00000000; // 
         11'h2d6: data <= 8'b00000000; // 
         11'h2d7: data <= 8'b01111110; //  ******
         11'h2d8: data <= 8'b00000000; // 
         11'h2d9: data <= 8'b00000000; // 
         11'h2da: data <= 8'b00000000; // 
         11'h2db: data <= 8'b00000000; // 
         11'h2dc: data <= 8'b00000000; // 
         11'h2dd: data <= 8'b00000000; // 
         11'h2de: data <= 8'b00000000; // 
         11'h2df: data <= 8'b00000000; // 
			//code x2f
         11'h2f0: data <= 8'b00000000; // 
         11'h2f1: data <= 8'b00000000; // 
         11'h2f2: data <= 8'b00000000; // 
         11'h2f3: data <= 8'b00000000; // 
         11'h2f4: data <= 8'b00000010; //       *
         11'h2f5: data <= 8'b00000110; //      **
         11'h2f6: data <= 8'b00001100; //     **
         11'h2f7: data <= 8'b00011000; //    **
         11'h2f8: data <= 8'b00110000; //   **
         11'h2f9: data <= 8'b01100000; //  **
         11'h2fa: data <= 8'b11000000; // **
         11'h2fb: data <= 8'b10000000; // *
         11'h2fc: data <= 8'b00000000; // 
         11'h2fd: data <= 8'b00000000; // 
         11'h2fe: data <= 8'b00000000; // 
         11'h2ff: data <= 8'b00000000; // 
         //code x30
         11'h300: data <= 8'b00000000; // 
         11'h301: data <= 8'b00000000; // 
         11'h302: data <= 8'b01111100; //  *****
         11'h303: data <= 8'b11000110; // **   **
         11'h304: data <= 8'b11000110; // **   **
         11'h305: data <= 8'b11001110; // **  ***
         11'h306: data <= 8'b11011110; // ** ****
         11'h307: data <= 8'b11110110; // **** **
         11'h308: data <= 8'b11100110; // ***  **
         11'h309: data <= 8'b11000110; // **   **
         11'h30a: data <= 8'b11000110; // **   **
         11'h30b: data <= 8'b01111100; //  *****
         11'h30c: data <= 8'b00000000; // 
         11'h30d: data <= 8'b00000000; // 
         11'h30e: data <= 8'b00000000; // 
         11'h30f: data <= 8'b00000000; // 
         //code x31
         11'h310: data <= 8'b00000000; // 
         11'h311: data <= 8'b00000000; // 
         11'h312: data <= 8'b00011000; // 
         11'h313: data <= 8'b00111000; // 
         11'h314: data <= 8'b01111000; //    **
         11'h315: data <= 8'b00011000; //   ***
         11'h316: data <= 8'b00011000; //  ****
         11'h317: data <= 8'b00011000; //    **
         11'h318: data <= 8'b00011000; //    **
         11'h319: data <= 8'b00011000; //    **
         11'h31a: data <= 8'b00011000; //    **
         11'h31b: data <= 8'b01111110; //    **
         11'h31c: data <= 8'b00000000; //    **
         11'h31d: data <= 8'b00000000; //  ******
         11'h31e: data <= 8'b00000000; // 
         11'h31f: data <= 8'b00000000; // 
         //code x32
         11'h320: data <= 8'b00000000; // 
         11'h321: data <= 8'b00000000; // 
         11'h322: data <= 8'b01111100; //  *****
         11'h323: data <= 8'b11000110; // **   **
         11'h324: data <= 8'b00000110; //      **
         11'h325: data <= 8'b00001100; //     **
         11'h326: data <= 8'b00011000; //    **
         11'h327: data <= 8'b00110000; //   **
         11'h328: data <= 8'b01100000; //  **
         11'h329: data <= 8'b11000000; // **
         11'h32a: data <= 8'b11000110; // **   **
         11'h32b: data <= 8'b11111110; // *******
         11'h32c: data <= 8'b00000000; // 
         11'h32d: data <= 8'b00000000; // 
         11'h32e: data <= 8'b00000000; // 
         11'h32f: data <= 8'b00000000; // 
         //code x33
         11'h330: data <= 8'b00000000; // 
         11'h331: data <= 8'b00000000; // 
         11'h332: data <= 8'b01111100; //  *****
         11'h333: data <= 8'b11000110; // **   **
         11'h334: data <= 8'b00000110; //      **
         11'h335: data <= 8'b00000110; //      **
         11'h336: data <= 8'b00111100; //   ****
         11'h337: data <= 8'b00000110; //      **
         11'h338: data <= 8'b00000110; //      **
         11'h339: data <= 8'b00000110; //      **
         11'h33a: data <= 8'b11000110; // **   **
         11'h33b: data <= 8'b01111100; //  *****
         11'h33c: data <= 8'b00000000; // 
         11'h33d: data <= 8'b00000000; // 
         11'h33e: data <= 8'b00000000; // 
         11'h33f: data <= 8'b00000000; // 
         //code x34
         11'h340: data <= 8'b00000000; // 
         11'h341: data <= 8'b00000000; // 
         11'h342: data <= 8'b00001100; //     **
         11'h343: data <= 8'b00011100; //    ***
         11'h344: data <= 8'b00111100; //   ****
         11'h345: data <= 8'b01101100; //  ** **
         11'h346: data <= 8'b11001100; // **  **
         11'h347: data <= 8'b11111110; // *******
         11'h348: data <= 8'b00001100; //     **
         11'h349: data <= 8'b00001100; //     **
         11'h34a: data <= 8'b00001100; //     **
         11'h34b: data <= 8'b00011110; //    ****
         11'h34c: data <= 8'b00000000; // 
         11'h34d: data <= 8'b00000000; // 
         11'h34e: data <= 8'b00000000; // 
         11'h34f: data <= 8'b00000000; // 
         //code x35
         11'h350: data <= 8'b00000000; // 
         11'h351: data <= 8'b00000000; // 
         11'h352: data <= 8'b11111110; // *******
         11'h353: data <= 8'b11000000; // **
         11'h354: data <= 8'b11000000; // **
         11'h355: data <= 8'b11000000; // **
         11'h356: data <= 8'b11111100; // ******
         11'h357: data <= 8'b00000110; //      **
         11'h358: data <= 8'b00000110; //      **
         11'h359: data <= 8'b00000110; //      **
         11'h35a: data <= 8'b11000110; // **   **
         11'h35b: data <= 8'b01111100; //  *****
         11'h35c: data <= 8'b00000000; // 
         11'h35d: data <= 8'b00000000; // 
         11'h35e: data <= 8'b00000000; // 
         11'h35f: data <= 8'b00000000; // 
         //code x36
         11'h360: data <= 8'b00000000; // 
         11'h361: data <= 8'b00000000; // 
         11'h362: data <= 8'b00111000; //   ***
         11'h363: data <= 8'b01100000; //  **
         11'h364: data <= 8'b11000000; // **
         11'h365: data <= 8'b11000000; // **
         11'h366: data <= 8'b11111100; // ******
         11'h367: data <= 8'b11000110; // **   **
         11'h368: data <= 8'b11000110; // **   **
         11'h369: data <= 8'b11000110; // **   **
         11'h36a: data <= 8'b11000110; // **   **
         11'h36b: data <= 8'b01111100; //  *****
         11'h36c: data <= 8'b00000000; // 
         11'h36d: data <= 8'b00000000; // 
         11'h36e: data <= 8'b00000000; // 
         11'h36f: data <= 8'b00000000; // 
         //code x37
         11'h370: data <= 8'b00000000; // 
         11'h371: data <= 8'b00000000; // 
         11'h372: data <= 8'b11111110; // *******
         11'h373: data <= 8'b11000110; // **   **
         11'h374: data <= 8'b00000110; //      **
         11'h375: data <= 8'b00000110; //      **
         11'h376: data <= 8'b00001100; //     **
         11'h377: data <= 8'b00011000; //    **
         11'h378: data <= 8'b00110000; //   **
         11'h379: data <= 8'b00110000; //   **
         11'h37a: data <= 8'b00110000; //   **
         11'h37b: data <= 8'b00110000; //   **
         11'h37c: data <= 8'b00000000; // 
         11'h37d: data <= 8'b00000000; // 
         11'h37e: data <= 8'b00000000; // 
         11'h37f: data <= 8'b00000000; // 
         //code x38
         11'h380: data <= 8'b00000000; // 
         11'h381: data <= 8'b00000000; // 
         11'h382: data <= 8'b01111100; //  *****
         11'h383: data <= 8'b11000110; // **   **
         11'h384: data <= 8'b11000110; // **   **
         11'h385: data <= 8'b11000110; // **   **
         11'h386: data <= 8'b01111100; //  *****
         11'h387: data <= 8'b11000110; // **   **
         11'h388: data <= 8'b11000110; // **   **
         11'h389: data <= 8'b11000110; // **   **
         11'h38a: data <= 8'b11000110; // **   **
         11'h38b: data <= 8'b01111100; //  *****
         11'h38c: data <= 8'b00000000; // 
         11'h38d: data <= 8'b00000000; // 
         11'h38e: data <= 8'b00000000; // 
         11'h38f: data <= 8'b00000000; // 
         //code x39
         11'h390: data <= 8'b00000000; // 
         11'h391: data <= 8'b00000000; // 
         11'h392: data <= 8'b01111100; //  *****
         11'h393: data <= 8'b11000110; // **   **
         11'h394: data <= 8'b11000110; // **   **
         11'h395: data <= 8'b11000110; // **   **
         11'h396: data <= 8'b01111110; //  ******
         11'h397: data <= 8'b00000110; //      **
         11'h398: data <= 8'b00000110; //      **
         11'h399: data <= 8'b00000110; //      **
         11'h39a: data <= 8'b00001100; //     **
         11'h39b: data <= 8'b01111000; //  ****
         11'h39c: data <= 8'b00000000; // 
         11'h39d: data <= 8'b00000000; // 
         11'h39e: data <= 8'b00000000; // 
         11'h39f: data <= 8'b00000000; // 
 endcase  
 
 
 always@*
	data_reg <= data;
 
   	       
endmodule